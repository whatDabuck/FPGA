module modulename #
// (

// )
(
    input a,b,
    output c
);
    reg a_tmp;
    reg b_tmp;

endmodule
module modulename #
// (

// )
(
    input a,b,
    output c
);



endmodule
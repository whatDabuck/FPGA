module modulename #
(

)
(
    ports
);
    
endmodule